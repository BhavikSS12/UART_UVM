// UART Corner Case Test
// File: tb/tests/uart_corner_test.sv

class uart_corner_test extends uart_base_test;
    
    `uvm_component_utils(uart_corner_test)
    
    function new(string name = "uart_corner_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction
    
    virtual task run_phase(uvm_phase phase);
        uart_corner_sequence seq;
        
        phase.raise_objection(this);
        
        super.run_phase(phase);
        
        `uvm_info(get_type_name(), "============================================", UVM_LOW)
        `uvm_info(get_type_name(), "  Starting Corner Case Test", UVM_LOW)
        `uvm_info(get_type_name(), "  Values: 0x00, 0xFF, 0xAA, 0x55, 0x0F, 0xF0", UVM_LOW)
        `uvm_info(get_type_name(), "============================================", UVM_LOW)
        
        seq = uart_corner_sequence::type_id::create("seq");
        seq.start(env.agent.sequencer);
        
        #5000;
        
        `uvm_info(get_type_name(), "Corner case test completed", UVM_LOW)
        
        phase.drop_objection(this);
    endtask
    
endclass